////////////////////////////////////////////////////////////////////////////////
// Type definitions
////////////////////////////////////////////////////////////////////////////////
`define E1__zero 2'h0
`define E1__first 2'h1
`define E1__second 2'h2
`define E1__third 2'h3





////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [14:0] in_a,
	output logic [1:0] out_a,
	output logic [14:0] out_b
);

	assign out_a = in_a;
	assign out_b = out_a;

endmodule


