////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [4:0] i,
	input logic [4:0] s,
	output logic o
);

	assign o = 
		(s[0] ? i[0] : 1'b0) | 
		(s[1] ? i[1] : 1'b0) | 
		(s[2] ? i[2] : 1'b0) | 
		(s[3] ? i[3] : 1'b0) | 
		(s[4] ? i[4] : 1'b0) ;

endmodule


