////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	output logic signed [4:0] out_a,
	input logic signed [2:0] in_a,
	input logic signed [2:0] in_b
);

	logic signed [3:0] u_output_port;

	assign out_a = u_output_port;

	DecoratorModule u (
		.output_port(u_output_port),
		.a(in_a),
		.b(in_b)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// DecoratorModule
////////////////////////////////////////////////////////////////////////////////
module DecoratorModule (
	output logic signed [3:0] output_port,
	input logic signed [2:0] a,
	input logic signed [2:0] b
);

	assign output_port = a + b;

endmodule


