////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [6:0] a_top,
	output logic [6:0] o_top,
	output logic [7:0] o2_top
);

	assign o2_top = 7'h7b;

	Sub u (
		.a_sub(o2_top)
	);

	assign o_top = a_top;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Sub
////////////////////////////////////////////////////////////////////////////////
module Sub (
	input logic [6:0] a_sub,
	output logic [7:0] o_sub
);

	assign o_sub = a_sub;
endmodule


