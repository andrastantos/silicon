////////////////////////////////////////////////////////////////////////////////
// Outer
////////////////////////////////////////////////////////////////////////////////
module Outer (
);

	logic wire2;
	logic wire1;

	Inner1 inner1 (
		.inner1_in(1'hx),
		.inner1_out1(wire1),
		.inner1_out2(wire2)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner1
////////////////////////////////////////////////////////////////////////////////
module Inner1 (
	input logic inner1_in,
	output logic inner1_out1,
	output logic inner1_out2
);

	assign inner1_out2 = inner1_out1;

	Inner2 inner2 (
		.inner2_out(inner1_out1)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner2
////////////////////////////////////////////////////////////////////////////////
module Inner2 (
	output logic inner2_out
);

	assign inner2_out = 1'h1;

endmodule


