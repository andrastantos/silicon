////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	input logic [7:0] in_a,
	output logic [7:0] out_h
);

	Parity u (
		.input_port(in_a),
		.output_port(out_h)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Parity
////////////////////////////////////////////////////////////////////////////////
module Parity (
	input logic [7:0] input_port,
	output logic output_port
);

	assign output_port = 1'hx;
endmodule


