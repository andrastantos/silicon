////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [31:0] i,
	input logic [4:0] s,
	output logic o
);

	always @(*) begin
		unique case (s)
			5'd0: o = i[0];
			5'd1: o = i[1];
			5'd2: o = i[2];
			5'd3: o = i[3];
			5'd4: o = i[4];
			5'd5: o = i[5];
			5'd6: o = i[6];
			5'd7: o = i[7];
			5'd8: o = i[8];
			5'd9: o = i[9];
			5'd10: o = i[10];
			5'd11: o = i[11];
			5'd12: o = i[12];
			5'd13: o = i[13];
			5'd14: o = i[14];
			5'd15: o = i[15];
			5'd16: o = i[16];
			5'd17: o = i[17];
			5'd18: o = i[18];
			5'd19: o = i[19];
			5'd20: o = i[20];
			5'd21: o = i[21];
			5'd22: o = i[22];
			5'd23: o = i[23];
			5'd24: o = i[24];
			5'd25: o = i[25];
			5'd26: o = i[26];
			5'd27: o = i[27];
			5'd28: o = i[28];
			5'd29: o = i[29];
			5'd30: o = i[30];
			5'd31: o = i[31];
			default: o = 1'hx;
		endcase
	end

endmodule


