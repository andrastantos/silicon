////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [7:0] in1,
	output logic [7:0] out1,
	input logic latch,
	input logic rst
);

	always_comb if (rst) out1 = 8'h0; else if (latch == 0) out1 = in1;

endmodule


