////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [7:0] in1,
	output logic [9:0] outp
);

	assign outp = { in1 + 8'h9 + 9'b0, 1'b0 };

endmodule


