////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic clk,
	input logic rst
);

	logic [7:0] p_outp_fwd;

	Producer p (
		.clk(clk),
		.rst(rst),
		.outp_fwd(p_outp_fwd)
	);

	Consumer c (
		.clk(clk),
		.rst(rst),
		.inp_fwd(p_outp_fwd)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Consumer
////////////////////////////////////////////////////////////////////////////////
module Consumer (
	input logic clk,
	input logic rst,
	input logic [7:0] inp_fwd
);

	logic [7:0] x;

	always_ff @(posedge clk) x <= rst ? 8'h0 : inp_fwd;

endmodule


////////////////////////////////////////////////////////////////////////////////
// Producer
////////////////////////////////////////////////////////////////////////////////
module Producer (
	input logic clk,
	input logic rst,
	output logic [7:0] outp_fwd
);

	logic [7:0] x;

	always_ff @(posedge clk) x <= rst ? 8'h0 : 8'(x + 1'h1 + 9'b0);

	assign outp_fwd = x;
endmodule


