////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic uout11,
	input logic uin1,
	input logic uin2
);

	logic u_output_port;

	assign uout11 = u_output_port[0];

	assign u_output_port = uin1 | uin2;
endmodule


