////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic in_1,
	output logic out_1
);

	logic out_1_1;

	assign out_1 = in_1;
	assign out_1_1 = in_1;
endmodule


