////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	output logic [7:0] out_1,
	output logic [7:0] out_1b,
	output logic [7:0] out_2
);

	assign out_1 = 8'hf;
	assign out_1b = 8'hf;

	assign out_2 = 8'hx;
endmodule


