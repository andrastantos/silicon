////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic in_1,
	input logic in_2,
	output logic out_1
);

	logic A_out_a;

	and_gate A (
		.in_a(1'hx),
		.in_b(1'hx),
		.out_a(A_out_a)
	);

	assign out_1 = 1'hx;
endmodule


////////////////////////////////////////////////////////////////////////////////
// and_gate
////////////////////////////////////////////////////////////////////////////////
module and_gate (
	input logic in_a,
	input logic in_b,
	output logic out_a
);
	assign out_a = in_a & in_b;
endmodule





