////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [7:0] o,
	input logic [3:0] i
);

	logic [3:0] top_if_rev;
	logic [7:0] top_if_fwd;

	mod mmm (
		.mod_out_fwd(top_if_fwd),
		.mod_out_rev(i)
	);

	assign top_if_rev = i;
	assign o = top_if_fwd;
endmodule


////////////////////////////////////////////////////////////////////////////////
// mod
////////////////////////////////////////////////////////////////////////////////
module mod (
	output logic [7:0] mod_out_fwd,
	input logic [3:0] mod_out_rev
);

	logic [7:0] x;

	assign x = 6'h2a & mod_out_rev;

	assign mod_out_fwd = x;
endmodule


