////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input E1 in_a,
	output E1 out_a
);

	assign out_a = first & in_a;

endmodule


