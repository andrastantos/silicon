////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [4:0] out1,
	input logic [1:0] in1
);

	assign out1 = {in1, 3'(in1)};

endmodule


