////////////////////////////////////////////////////////////////////////////////
// Outer
////////////////////////////////////////////////////////////////////////////////
module Outer (
);

	logic loopback;
	logic u_inner_out;

	assign loopback = u_inner_out;

	Inner u (
		.inner_in(loopback),
		.inner_out(u_inner_out)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner
////////////////////////////////////////////////////////////////////////////////
module Inner (
	input logic inner_in,
	output logic inner_out
);

	assign inner_out = 1'h1;

endmodule


