////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [1:0] sout1,
	input logic [1:0] uin1,
	input logic clk
);

	always_ff @(posedge clk) sout1 <= uin1;

endmodule


