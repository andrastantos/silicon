////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
);

	logic [31:0] c2bus_data_out;
	logic [31:0] c1bus_data_out;

	Procuder producer (
		.fetch_data_out(c1bus_data_out),

		.mem_data_out(c2bus_data_out)
	);

	Consumer1 consumer1 (
		.bus_if_data_out(c1bus_data_out)
	);

	Consumer2 consumer2 (
		.bus_if_data_out(c2bus_data_out)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Consumer2
////////////////////////////////////////////////////////////////////////////////
module Consumer2 (
	input logic [31:0] bus_if_data_out
);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Consumer1
////////////////////////////////////////////////////////////////////////////////
module Consumer1 (
	input logic [31:0] bus_if_data_out
);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Procuder
////////////////////////////////////////////////////////////////////////////////
module Procuder (
	output logic [31:0] fetch_data_out,
	output logic [31:0] mem_data_out
);

	logic [31:0] data_out;

	assign data_out = 1'h1;
	assign fetch_data_out = data_out;

	assign mem_data_out = data_out;
endmodule


