////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [1:0] uout1,
	output logic [1:0] uout2,
	input logic [1:0] uin1
);

	assign uout1 = {uin1[1], uin1[0]};

	assign uout2 = 2'hx;
endmodule


