////////////////////////////////////////////////////////////////////////////////
// Outer
////////////////////////////////////////////////////////////////////////////////
module Outer (
);

	logic inner1_inner1_out;
	logic inner2_inner2_out;

	Inner2 inner2 (
		.inner2_in(inner1_inner1_out),
		.inner2_out(inner2_inner2_out)
	);

	Inner1 inner1 (
		.inner1_in(inner2_inner2_out),
		.inner1_out(inner1_inner1_out)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner1
////////////////////////////////////////////////////////////////////////////////
module Inner1 (
	input logic inner1_in,
	output logic inner1_out
);

	assign inner1_out = 1'hx;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner2
////////////////////////////////////////////////////////////////////////////////
module Inner2 (
	input logic inner2_in,
	output logic inner2_out
);

	assign inner2_out = inner2_in;

endmodule


