////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic signed [7:0] input,
	output logic signed [7:0] output1,
	output logic signed [7:0] output2
);

	assign output2 = 1'h0;

	assign output1 = input;
endmodule


