////////////////////////////////////////////////////////////////////////////////
// Outer
////////////////////////////////////////////////////////////////////////////////
module Outer (
	input logic outer_in,
	output logic outer_out
);

	Inner u (
		.inner_in(outer_in),
		.inner_out(outer_out)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner
////////////////////////////////////////////////////////////////////////////////
module Inner (
	input logic inner_in,
	output logic inner_out
);

	assign inner_out = inner_in;

endmodule


