////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	output logic [4:0] out_a,
	output logic [4:0] out_b,
	input logic [2:0] in_a,
	input logic [2:0] in_b
);

	DecoratorModule u (
		.output_port(out_a),
		.a(in_a)
	);

	DecoratorModule_2 u3 (
		.output_port(out_b),
		.a(in_a[2:0]),
		.b(in_b[1])
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// DecoratorModule_2
////////////////////////////////////////////////////////////////////////////////
module DecoratorModule_2 (
	output logic [3:0] output_port,
	input logic [2:0] a,
	input logic b
);

	assign output_port = a + b;

endmodule


////////////////////////////////////////////////////////////////////////////////
// DecoratorModule
////////////////////////////////////////////////////////////////////////////////
module DecoratorModule (
	output logic output_port,
	input logic [2:0] a
);

	assign output_port = a[0];

endmodule


