////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [1:0] a,
	input logic [2:0] b,
	input logic [3:0] c,
	input logic [4:0] d,
	output logic [7:0] o
);

	assign o = {c[3], b, a[0], 3'(a)};

endmodule


