////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic signed [7:0] input_port,
	output logic signed [7:0] output_port
);

	assign output_port = 8'hx;
endmodule


