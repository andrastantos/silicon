////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic signed [4:0] out_a,
	input logic signed in_a,
	input logic signed in_b
);

	assign out_a = $signed({in_a & in_b, 2'(1'h1), 2'(1'h0)});

endmodule


