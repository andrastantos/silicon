////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [7:0] a,
	output logic [7:0] o,
	output logic [7:0] o2
);

	Sub u (
		.o(o2)
	);

	assign o = a;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Sub
////////////////////////////////////////////////////////////////////////////////
module Sub (
	output logic [7:0] o
);

	logic [7:0] a;

	assign o = a;
	assign a = 123;
endmodule


