////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic signed [7:0] input,
	output logic signed [7:0] output
);

	assign output = 8'x;
endmodule


