////////////////////////////////////////////////////////////////////////////////
// Outer
////////////////////////////////////////////////////////////////////////////////
module Outer (
);

	logic u1_output_port;
	logic loopback;

	Inner u (
		.inner_in(u1_output_port),
		.inner_out(loopback)
	);

	assign u1_output_port = loopback;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Inner
////////////////////////////////////////////////////////////////////////////////
module Inner (
	input logic inner_in,
	output logic inner_out
);

	assign inner_out = 1'h1;

endmodule


