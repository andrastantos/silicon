////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	input logic [7:0] in_a,
	output logic [7:0] out_h
);

	logic u_output;

	assign out_h = u_output;

	Parity u (
		.input(in_a),
		.output(u_output)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Parity
////////////////////////////////////////////////////////////////////////////////
module Parity (
	input logic [7:0] input,
	output logic output
);

endmodule


