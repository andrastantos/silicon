////////////////////////////////////////////////////////////////////////////////
// Type definitions
////////////////////////////////////////////////////////////////////////////////
typedef enum logic [1:0] {
	first=1,
	second=2,
	third=3
} E1;




////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input E1 in_a,
	output E1 out_a
);

	assign out_a = in_a;
endmodule


