////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	input logic [7:0] in_a,
	output logic [7:0] out_1,
	output logic [7:0] out_2,
	output logic [7:0] out_3
);

	Parity u (
		.input(in_a),
		.output(out_1)
	);

	Parity u1 (
		.input(in_a),
		.output(out_2)
	);

	assign out_3 = 8'bX;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Parity
////////////////////////////////////////////////////////////////////////////////
module Parity (
	input logic [7:0] input,
	output logic output
);

	assign output = input[0];

endmodule


