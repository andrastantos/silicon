////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic top_in1,
	input logic top_in2,
	output logic top_out
);

	logic yyy;
	logic xxx;

	assign xxx = top_in1 & top_in2;

	assign top_out = xxx;
	assign yyy = xxx;
endmodule


