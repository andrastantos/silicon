////////////////////////////////////////////////////////////////////////////////
// test_module
////////////////////////////////////////////////////////////////////////////////
module test_module (
	input logic [1:0] data_in
);

endmodule


