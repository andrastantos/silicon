////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	output logic [4:0] out_a,
	input logic in_c
);

	logic [3:0] x;

	assign x = out_a[3:0];
	assign out_a = {1'h1, 4'(in_c)};

endmodule


