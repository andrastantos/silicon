////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic top_in_bwd,
	input logic [1:0] top_in_fwd
);

	logic [1:0] top_w_fwd;
	logic top_w_bwd;

	assign top_w_bwd = 1'h1;

	assign top_w_fwd = top_in_fwd;
	assign top_in_bwd = top_w_bwd;
endmodule


