////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [6:0] a_top,
	output logic [6:0] o_top,
	output logic [7:0] o2_top
);

	logic [6:0] u3_output_port;

	assign o_top = a_top;

	Sub u (
		.a_sub(u3_output_port),
		.o_sub(o2_top)
	);

	assign u3_output_port = 7'h7b;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Sub
////////////////////////////////////////////////////////////////////////////////
module Sub (
	input logic [6:0] a_sub,
	output logic [7:0] o_sub
);

	assign o_sub = a_sub;

endmodule


