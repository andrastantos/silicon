////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic top_in1,
	input logic top_in2,
	output logic top_out
);

	logic xxx;
	logic yyy;

	assign yyy = top_in1 & top_in2;

	assign top_out = yyy;
	assign xxx = yyy;
endmodule


