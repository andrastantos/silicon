////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic uout1,
	output logic uout2,
	input logic [1:0] uin1
);

	logic x;

	assign x = uin1[0];
	assign uout1 = uin1[1];

	assign uout2 = x;
endmodule


