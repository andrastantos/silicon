////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [3:0] in1,
	input logic [3:0] in2,
	input logic sel,
	output logic [3:0] out1
);

	assign out1 = sel ? in2 : in1;

endmodule


