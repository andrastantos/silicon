////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [7:0] i1,
	input logic i2,
	output logic o
);

	assign o = i2 & i1 == 6'h2a;

endmodule


