////////////////////////////////////////////////////////////////////////////////
// Type definitions
////////////////////////////////////////////////////////////////////////////////
`define E1__first 2'h1
`define E1__second 2'h2
`define E1__third 2'h3





////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [1:0] in_a,
	output logic [1:0] out_a
);

	assign out_a = `E1__first & in_a;

endmodule


