////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic in_a,
	output logic out_a
);

	and_gate A (
		.in_a(in_a),
		.in_b(in_a),
		.out_a(out_a)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// and_gate
////////////////////////////////////////////////////////////////////////////////
module and_gate (
	input logic in_a,
	input logic in_b,
	output logic out_a
);

	assign out_a = 1'hx;
endmodule


