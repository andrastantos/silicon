////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic [3:0] i,
	output logic [5:0] o
);

	logic [3:0] top_if_rev;

	mod mmm (
		.mod_out_rev(i),

		.x(o)
	);

	assign top_if_rev = i;
endmodule


////////////////////////////////////////////////////////////////////////////////
// mod
////////////////////////////////////////////////////////////////////////////////
module mod (
	input logic [3:0] mod_out_rev,
	output logic [5:0] x
);

	assign x = 6'h2a & mod_out_rev;

endmodule


