////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input E1 in_a,
	output logic [1:0] out_a
);

	assign out_a = first & in_a;

endmodule


