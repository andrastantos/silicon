////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic [7:0] i1,
	output logic [4:0] o
);

	assign o = i1[3:0];

endmodule


