////////////////////////////////////////////////////////////////////////////////
// Top
////////////////////////////////////////////////////////////////////////////////
module Top (
	input logic signed [7:0] in1,
	input logic [7:0] in2,
	output logic signed [9:0] outp
);

	assign outp = { in1, 1'b0 } + in2 + 10'b0 >>> 1;

endmodule


