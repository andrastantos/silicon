////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [31:0] push_data
);

	assign push_data = 2'h3;

endmodule


