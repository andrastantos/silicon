////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	input logic [7:0] in_a,
	output logic [7:0] out_h
);

	logic u_output_port;

	assign out_h = u_output_port;

	Parity u (
		.input_port(in_a),
		.output_port(u_output_port)
	);

endmodule


////////////////////////////////////////////////////////////////////////////////
// Parity
////////////////////////////////////////////////////////////////////////////////
module Parity (
	input logic [7:0] input_port,
	output logic output_port
);

	assign output_port = 1'x;
endmodule


