////////////////////////////////////////////////////////////////////////////////
// Test
////////////////////////////////////////////////////////////////////////////////
module Test (
	input logic [7:0] in_a,
	output logic [7:0] out_1,
	output logic [7:0] out_2,
	output logic [7:0] out_3
);

	Parity u (
		.input_port(in_a),
		.output_port(out_1)
	);

	Parity u1 (
		.input_port(in_a),
		.output_port(out_2)
	);

	assign out_3 = 8'x;
endmodule


////////////////////////////////////////////////////////////////////////////////
// Parity
////////////////////////////////////////////////////////////////////////////////
module Parity (
	input logic [7:0] input_port,
	output logic output_port
);

	assign output_port = input_port[0];

endmodule


