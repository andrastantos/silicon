////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic uout11,
	input logic uin1,
	input logic uin2
);

	assign uout11 = (uin1 | uin2)[0];

endmodule


