////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	output logic [7:0] out_a,
	input logic [7:0] in_a
);

	assign out_a = {7'(1'h1), in_a[0]};

endmodule


