////////////////////////////////////////////////////////////////////////////////
// top
////////////////////////////////////////////////////////////////////////////////
module top (
	input logic top_port,
	output logic top_out
);

	assign top_out = top_port;

endmodule


